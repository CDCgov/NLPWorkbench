Clinical History||(?:^[\t ]*CLINICAL HISTORY):?\r?\n
Family History||(?:^[\t ]*FAMILY HISTORY):?\r?\n
History of Present Illness||(?:^[\t ]*(?:(?:HISTORY OF PAST ILLNESS)|(?:PAST MEDICAL HISTORY))):?\r?\n
History of Present Illness||(?:^[\t ]*(?:HISTORY OF PRESENT ILLNESS| history of physical illness,history of present illness,history of the present illness)):?\r?\n
